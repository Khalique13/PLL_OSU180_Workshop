* SPICE3 file created from std_cells.ext - technology: scmos

.option scale=0.1u

M1000 w_632_550# a_660_506# a_655_556# w_632_550# pfet w=11 l=2
+  ad=0 pd=0 as=0 ps=0
M1001 a_655_556# a_648_496# w_632_550# w_632_550# pfet w=11 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 a_563_489# a_556_520# a_556_488# a_556_488# nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_777_556# a_795_526# a_788_484# a_556_488# nfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_788_484# a_782_521# a_777_484# a_556_488# nfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 a_777_484# a_774_532# a_556_488# a_556_488# nfet w=9 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 a_777_556# a_795_526# w_760_550# w_760_550# pfet w=11 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 a_655_556# a_660_506# a_655_487# a_556_488# nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 w_760_550# a_782_521# a_777_556# w_760_550# pfet w=11 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a_777_556# a_774_532# w_760_550# w_760_550# pfet w=11 l=2
+  ad=0 pd=0 as=0 ps=0
M1010 a_563_489# a_556_520# w_550_550# w_550_550# pfet w=11 l=2
+  ad=0 pd=0 as=0 ps=0
M1011 a_655_487# a_648_496# a_556_488# a_556_488# nfet w=6 l=2
+  ad=0 pd=0 as=0 ps=0
C0 a_782_521# a_777_556# 0.01fF
C1 a_782_521# w_760_550# 0.07fF
C2 a_774_532# a_795_526# 0.01fF
C3 w_550_550# a_563_489# 0.18fF
C4 a_782_521# a_774_532# 0.08fF
C5 a_777_556# w_760_550# 0.33fF
C6 a_648_496# a_660_506# 0.13fF
C7 a_655_556# a_660_506# 0.13fF
C8 a_563_489# a_556_520# 0.05fF
C9 a_782_521# a_795_526# 0.02fF
C10 a_648_496# w_632_550# 0.07fF
C11 a_655_556# w_632_550# 0.21fF
C12 a_660_506# w_632_550# 0.07fF
C13 a_774_532# w_760_550# 0.07fF
C14 w_550_550# a_556_520# 0.07fF
C15 a_795_526# a_777_556# 0.08fF
C16 a_795_526# w_760_550# 0.07fF
C17 a_777_556# a_556_488# 0.35fF
C18 a_655_556# a_556_488# 0.27fF
C19 a_563_489# a_556_488# 0.28fF
C20 a_795_526# a_556_488# 0.49fF
C21 a_782_521# a_556_488# 0.53fF
C22 a_774_532# a_556_488# 0.50fF
C23 a_660_506# a_556_488# 0.52fF
C24 a_648_496# a_556_488# 0.56fF
C25 a_556_520# a_556_488# 0.49fF
C26 w_760_550# a_556_488# 1.80fF
C27 w_632_550# a_556_488# 1.83fF
C28 w_550_550# a_556_488# 0.98fF
