* SPICE3 file created from inv.ext - technology: scmos

.option scale=0.1u

M1000 out in vdd vdd pfet w=8 l=2
+  ad=0 pd=0 as=0 ps=0
M1001 out in gnd gnd nfet w=3 l=2
+  ad=0 pd=0 as=0 ps=0
C0 in out 0.05fF
C1 out vdd 0.12fF
C2 in vdd 0.09fF
C3 out gnd 0.28fF
C4 in gnd 0.49fF
C5 vdd gnd 0.98fF
